
`timescale 1 ns / 1 ps

module s_axi_stream(/*AUTOARG*/
   // Outputs
   tready, buf_we, buf_wdata,
   // Inputs
   clk, xrst, tvalid, tdata, tstrb, tlast, buf_isfull
   );
`include "parameters.vh"

  parameter WORDS = 2 ** BUFSIZE;

  localparam  S_IDLE  = 'd0,
              S_WRITE = 'd1;

  /*AUTOINPUT*/
  input                 clk;
  input                 xrst;
  input                 tvalid;
  input [DWIDTH-1:0]    tdata;
  input [DWIDTH/8-1:0]  tstrb;
  input                 tlast;
  input                 buf_isfull;

  /*AUTOOUTPUT*/
  output              tready;
  output              buf_we;
  output [DWIDTH-1:0] buf_wdata;

  /*AUTOWIRE*/
  wire s_write_end;

  /*AUTOREG*/
  reg r_state;
  reg r_tready;
  reg r_write_end;

//==========================================================
// core control
//==========================================================

  always @(posedge clk)
    if (!xrst)
      r_state <= S_IDLE;
    else
      case (r_state)
        S_IDLE:
          if (tvalid)
            r_state <= S_WRITE;

        S_WRITE:
          if (s_write_end)
            r_state <= S_IDLE;
      endcase

//==========================================================
// stream control
//==========================================================

  assign tready = r_tready;

  always @(posedge clk)
    if (!xrst)
      r_tready <= 0;
    else
      r_tready <= r_state == S_WRITE && !buf_isfull;

//==========================================================
// buffer control
//==========================================================

  assign s_write_end = r_write_end;

  assign buf_we    = tvalid && r_tready;
  assign buf_wdata = tdata;

  always @(posedge clk)
    if (!xrst)
      r_write_end <= 0;
    else
      if (!buf_isfull) begin
        if (buf_we)
          r_write_end <= 0;
        if (buf_isfull || tlast)
          r_write_end <= 1;
      end

endmodule

